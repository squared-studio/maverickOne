/*
Description
Author : S. M. Tahmeed Reza (https://github.com/tahmeedKENJI)
This file is part of squared-studio:maverickOne
Copyright (c) 2025 squared-studio
Licensed under the MIT License
See LICENSE file in the project root for full license information
*/

module priority_encoder_tb;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-IMPORTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // bring in the testbench essentials functions and macros
  `include "vip/tb_ess.sv"

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  localparam int NumWire = 16;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  typedef logic [NumWire-1:0] n_wire;
  typedef logic [$clog2(NumWire)-1:0] n_encode;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // generates static task start_clk_i with tHigh:4ns tLow:6ns
  `CREATE_CLK(clk_i, 4ns, 6ns)

  n_wire wire_in;
  n_encode index_o;
  logic index_valid_o;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-VARIABLES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  int pen_counter;
  bit priority_violation_flag;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  priority_encoder #(
      .NUM_WIRE(NumWire)
  ) u_pen1 (
      .wire_in,
      .index_o,
      .index_valid_o
  );

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  task automatic start_random_driver();
    fork
      forever begin
        @(posedge clk_i);
        wire_in <= $urandom;
        pen_counter++;
      end
    join_none
  endtask

  task automatic start_in_out_monitor();
    pen_counter = 0;
    priority_violation_flag = 0;
    fork
      forever begin
        logic valid;
        @(posedge clk_i);
        valid = |wire_in;

        if (valid === '1) begin
          if ((index_valid_o === valid) && (index_o === priority_idx())) begin
            pen_counter++;
          end else begin
            priority_violation_flag = 1;
            result_print(0, "Priority Encoding Failed");
            $finish;
          end
        end
      end
    join_none
  endtask

  function automatic integer priority_idx();
    for (integer i = 0; i < NumWire; i++) begin
      if (wire_in[i] === '1) return i;
    end
  endfunction

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-PROCEDURALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  initial begin  // main initial
    start_clk_i();
    start_random_driver();
    start_in_out_monitor();
    repeat (1000) @(posedge clk_i);
    result_print(!priority_violation_flag, "Priority Encoding");
    $finish;
  end

endmodule
