/*
The `branch_target_buffer` is designed to store and manage branch target addresses for a processor,
helping to predict the next instruction address in case of a branch or jump.
Author : Subhan Zawad Bihan (https://github.com/SubhanBihan)
This file is part of squared-studio:maverickOne
Copyright (c) 2025 squared-studio
Licensed under the MIT License
See LICENSE file in the project root for full license information
*/

`include "maverickOne_pkg.sv"

module branch_target_buffer #(
    parameter int NUM_BTBL = maverickOne_pkg::NUM_BTBL,  // Number of branch target buffer lines
    parameter int XLEN     = maverickOne_pkg::XLEN       // Integer register width
) (
    input logic clk_i,   // Clock input
    input logic arst_ni, // Asynchronous reset input

    input logic [XLEN-1:0] current_addr_i,  // Current address (EXEC) input
    input logic [XLEN-1:0] next_addr_i,     // Next address (EXEC) input
    input logic [XLEN-1:0] pc_i,            // Program counter (IF) input
    input logic            is_jump_i,       // Is jump/branch (IF) input

    output logic            match_found_o,   // Found match in buffer output
    output logic            update_table_o,  // Table update event output
    output logic [XLEN-1:0] next_pc_o        // Next program counter (in case of jump) output
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  typedef logic [XLEN-1:2] reduced_addr_t;  // Reduced address type (excluding last 2 bits)

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  ///////////////////////////////////////////////
  // REGISTERS
  ///////////////////////////////////////////////

  // Buffer to store current addresses
  reduced_addr_t current_addr_buffer[NUM_BTBL];
  // Buffer to store next addresses
  reduced_addr_t next_addr_buffer[NUM_BTBL];
  // Valid bits for buffer entries
  logic [NUM_BTBL-1:0] valid_buffer;
  // Counter for buffer entries
  logic [$clog2(NUM_BTBL)-1:0] buffer_counter;

  ///////////////////////////////////////////////
  // WIRES
  ///////////////////////////////////////////////

  // Write enable signals for buffer entries
  logic [NUM_BTBL-1:0] write_enable;

  // Flag to check if next address is not equal to current address + 4
  logic addr_mismatch;

  // Match signals for program counter and current address
  logic [NUM_BTBL-1:0] pc_addr_match;
  // Index of matching row in buffer
  logic [$clog2(NUM_BTBL)-1:0] match_index;
  // Index of empty row in buffer
  logic [$clog2(NUM_BTBL)-1:0] empty_index;
  // Index of row to write in buffer
  logic [$clog2(NUM_BTBL)-1:0] write_index;

  // Flag to indicate if an empty row is found
  logic empty_found;
  // Flag to indicate if a match is found
  logic match_found;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // Check for matches between program counter and current addresses in buffer
  for (genvar i = 0; i < NUM_BTBL; i++) begin : g_pc_addr_match
    always_comb pc_addr_match[i] = valid_buffer[i] & (pc_i == current_addr_buffer[i]);
  end

  // Output match_found signal if a match is found or table is updated
  always_comb match_found_o = match_found | update_table_o;

  // Output next program counter based on table update or buffer content
  always_comb next_pc_o = update_table_o ? next_addr_i : {next_addr_buffer[match_index], 2'b00};

  // Check if next address is not equal to current address + 4
  always_comb addr_mismatch = (current_addr_i + 4 != next_addr_i);

  // Update table if there is a jump and addresses do not match
  always_comb update_table_o = is_jump_i & (addr_mismatch ^ match_found);

  // Determine the row index to write in buffer
  always_comb
    write_index = addr_mismatch ? (empty_found ? empty_index : buffer_counter) : match_index;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // Instance of the demux module to generate write enable signals
  demux #(
      .NUM_ELEM  (NUM_BTBL),
      .ELEM_WIDTH(1)
  ) u_demux (
      .index_i(write_index),
      .data_i (update_table_o),
      .out_o  (write_enable)
  );

  // Instance of the encoder module to find matching row index
  encoder #(
      .NUM_WIRE(NUM_BTBL)
  ) pc_addr_match_find (
      .wire_in(pc_addr_match),
      .index_o(match_index),
      .index_valid_o(match_found)
  );

  // Instance of the priority encoder module to find empty row index
  priority_encoder #(
      .NUM_WIRE(NUM_BTBL)
  ) empty_row_find (
      .wire_in(~valid_buffer),
      .index_o(empty_index),
      .index_valid_o(empty_found)
  );

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // Sequential logic to update buffer entries
  for (genvar i = 0; i < NUM_BTBL; i++) begin : g_regs
    always @(posedge clk_i) begin
      if (write_enable[i]) begin
        current_addr_buffer[i] <= current_addr_i[XLEN-1:2];
      end
    end

    always @(posedge clk_i) begin
      if (write_enable[i]) begin
        next_addr_buffer[i] <= next_addr_i[XLEN-1:2];
      end
    end

    // Sequential logic to update valid bits for buffer entries
    always_ff @(posedge clk_i or negedge arst_ni) begin
      if (~arst_ni) begin
        valid_buffer[i] <= '0;
      end else if (write_enable[i]) begin
        valid_buffer[i] <= addr_mismatch;
      end
    end
  end

  // Sequential logic to update counter
  always_ff @(posedge clk_i or negedge arst_ni) begin
    if (~arst_ni) begin
      buffer_counter <= '0;
    end else begin
      if (~empty_found & is_jump_i) buffer_counter <= buffer_counter + 1;
    end
  end

endmodule
