/*
The maverickOne module is designed to interface with instruction and data caches in a RISC-V 64-bit
architecture. It handles memory requests, data transfers, and interrupt management, making it
essential for efficient processor operation. Here's a detailed description of its functionality:
- **Memory Requests**: Manages requests to instruction and data caches, ensuring proper data flow
  between the processor and memory.
- **Data Transfers**: Handles data transfers to and from the caches, including specifying the
  address and size of the data.
- **Interrupt Management**: Processes interrupt requests, determines the active interrupt, and
  acknowledges interrupts, ensuring timely and efficient interrupt handling.
Author : Foez Ahmed (https://github.com/foez-ahmed)
This file is part of DSInnovators:maverickOne
Copyright (c) 2024 DSInnovators
Licensed under the MIT License
See LICENSE file in the project root for full license information
*/

module maverickOne #(
    localparam int AW   = 64,  // Address width
    localparam int ICDW = 32,  // I-Cache data width
    localparam int DCDW = 64   // D-Cache data width
) (
    input logic arst_ni,  // Asynchronous reset, active low
    input logic clk_i,    // Clock input

    // I-Cache Interface
    output logic            icache_req_o,   // I-Cache request signal
    output logic [  AW-1:0] icache_addr_o,  // I-Cache address output
    input  logic [ICDW-1:0] icache_data_i,  // I-Cache data input
    input  logic            icache_gnt_i,   // I-Cache grant signal

    // D-Cache Interface
    output logic            dcache_req_o,   // D-Cache request signal
    output logic            dcache_wr_o,    // D-Cache write/read signal
    output logic [  AW-1:0] dcache_addr_o,  // D-Cache address output
    output logic [     1:0] dcache_size_o,  // D-Cache size output
    output logic [DCDW-1:0] dcache_data_o,  // D-Cache data output
    input  logic [DCDW-1:0] dcache_data_i,  // D-Cache data input
    input  logic            dcache_gnt_i,   // D-Cache grant signal

    // Interrupt Interface
    input  logic [31:0] int_req_i,    // Interrupt request signals
    output logic [ 4:0] int_index_o,  // Interrupt index output
    output logic        int_ack_o     // Interrupt acknowledge signal
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS GENERATED
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INITIAL CHECKS
  //////////////////////////////////////////////////////////////////////////////////////////////////

endmodule
